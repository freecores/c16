library IEEE;
use IEEE.STD_LOGIC_1164.all;

package mem_content is

-- content of m_0_0
constant m_0_0_0 : BIT_VECTOR := X"3E5FFDDF2E8FF7FF56FFF56A97FFAB511FFEAD4066EFB555B5B6BB6A38000098";
constant m_0_0_1 : BIT_VECTOR := X"0A9A999AADED9BDB7E3C2C87F7FEACF6FFEEF6E567B7FF77B62B3E5FFDDF2E8B";
constant m_0_0_2 : BIT_VECTOR := X"A779CB7BD6BF6AA4B964EFAFC00786D5BB6EEA50AB24DB77C25B1A3DF1976DDD";
constant m_0_0_3 : BIT_VECTOR := X"9C9784DEA0DDC979FF93756424A1F89C979FF83752424B557F5FD7F5795E569D";
constant m_0_0_4 : BIT_VECTOR := X"C29BD98577B31415BD9062CF9ABC563B93B89C979FF93752424325E7FE4DD590";
constant m_0_0_5 : BIT_VECTOR := X"E2D627F5A9F6AD93BFAD85098577B30A6F6615DECC29BD98577B30A6F6615DEC";
constant m_0_0_6 : BIT_VECTOR := X"FC494DCADA963F4928E23FEF39FD9ABF7747C65D0AB43A1468556A569E5EB3F5";
constant m_0_0_7 : BIT_VECTOR := X"AEAB296639435AF7B5A739CEF79CFDED6F7E4B4EBDF95B528D6DDD9BB366EC55";
constant m_0_0_8 : BIT_VECTOR := X"15AA802B557C9444A294A1092C9253DF9FA51CE944962BA51CE944B3D2CE74A2";
constant m_0_0_9 : BIT_VECTOR := X"4656F56AF5AAD1AB7B323CD54923EDD8B55628CB91342F285BA4A26600920404";
constant m_0_0_A : BIT_VECTOR := X"000000000000000000000000000000000000000000000000000AA8BAB558C8AE";
constant m_0_0_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_1
constant m_0_1_0 : BIT_VECTOR := X"AA42949522A4D14B4C14B4C890A5A644429699012F2B49D9CFE23801D80001F8";
constant m_0_1_1 : BIT_VECTOR := X"E5AF0A8C6203045C2290E304D14A06AA14A4AA0C3510A5251021AA42949522A1";
constant m_0_1_2 : BIT_VECTOR := X"AD39DB5BD7BE90408B30ABE360003BFBA802AD2D7A9D4015E8D4870579D50055";
constant m_0_1_3 : BIT_VECTOR := X"6215726E91B42156F7D6D15BD89E4C62156F7C6D35392891CAD79CAD79CAD79D";
constant m_0_1_4 : BIT_VECTOR := X"13722C26A458519B22C509162809FCEE42AF62156F7D6D353928855BDF1B456F";
constant m_0_1_5 : BIT_VECTOR := X"58B5AB0DA5E97642AE5226F626A4584D48B09B91613722C26A4584D48B09B916";
constant m_0_1_6 : BIT_VECTOR := X"971E89A800E892E1D5AC1F9F2CA1A53F15F2B60FDF1F9FBF3F1F3E7EEDB58ED5";
constant m_0_1_7 : BIT_VECTOR := X"1C9C9EA011CB5AD694AF794A7394BDEFFB56F547B82F24BD1C0056AAB26AB614";
constant m_0_1_8 : BIT_VECTOR := X"2633004C665BEA2F467744E5D5CFA132E97A075E82E8857AB75E83C8BD03AF46";
constant m_0_1_9 : BIT_VECTOR := X"0119824165A34084C02040D19405253022204089820218401328840401203890";
constant m_0_1_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000014010048802126";
constant m_0_1_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_2
constant m_0_2_0 : BIT_VECTOR := X"922845C9119614230D4230D4CA11862228461A98A20721540C810CD09FFFFAD8";
constant m_0_2_1 : BIT_VECTOR := X"48C8A2008F10722681C38E7E1422DE41422E4132F24A117248D7902845C81117";
constant m_0_2_2 : BIT_VECTOR := X"128620A0280ED6E59B64873ADFFFE7602040704203890203121E2060C604080E";
constant m_0_2_3 : BIT_VECTOR := X"8898ED4A9534898DDA44D237225CE24898DDA44D27F6AA4421096B5AC4218D42";
constant m_0_2_4 : BIT_VECTOR := X"695906D2B20DB34B906BB7ECD9F6CB65121C8898DDA54D27F6AA2637695348DC";
constant m_0_2_5 : BIT_VECTOR := X"B6672C8EC0ED0D121D1AD2C8D2B20DA5641B4BC83697906D2F20DA5E41B4AC83";
constant m_0_2_6 : BIT_VECTOR := X"D6418DA011189ACA31B2F21327C846E4033DFE1CF9C339738652A70EDF6BFA41";
constant m_0_2_7 : BIT_VECTOR := X"05C78184970000002948429484295AD634FA0D58CFF6020350080E81D6A0772C";
constant m_0_2_8 : BIT_VECTOR := X"383C0070786C1A00D008C4A2314063C27B8613C1811AA38613C1A079C309E0C3";
constant m_0_2_9 : BIT_VECTOR := X"2A44F2EA8988BB2A788ABAC44FC298DD85972805093A0F28804472110192143C";
constant m_0_2_A : BIT_VECTOR := X"000000000000000000000000000000000000000000000000000B28D2365D4A94";
constant m_0_2_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_3
constant m_0_3_0 : BIT_VECTOR := X"2484441240011222EC222EC0011176840445DA10082A20110930004280000209";
constant m_0_3_1 : BIT_VECTOR := X"4808C465AA000643100BAB791222089C22209C2844A11104A00225844412C042";
constant m_0_3_2 : BIT_VECTOR := X"2B0A46908564D6E4A92F2A045FFFE5B14042A240088A02159244408540080854";
constant m_0_3_3 : BIT_VECTOR := X"A5EC444ABF355EC7DB7CD516695A7425EC7DB7CD5566B500D63485214A42918C";
constant m_0_3_4 : BIT_VECTOR := X"2542724A84E4952A272497A74AA24120BCA9A5EC7DB7CD5566BD7B1F6DF35459";
constant m_0_3_5 : BIT_VECTOR := X"0235888B704D24BCA89A4A9A4AC4E49589C92A1392542724A84E49509C92A139";
constant m_0_3_6 : BIT_VECTOR := X"404AD41010AFC8495B12E48BAA8800C915109710089020102041624FA1B02C91";
constant m_0_3_7 : BIT_VECTOR := X"C4AA8AF40836F79CC6318EF7BDE72948C65256888BC80215A808570A8A02B806";
constant m_0_3_8 : BIT_VECTOR := X"00C002018014AF856B156CB15F62BD22892B544AF8ADB12B544AF8A895EA256A";
constant m_0_3_9 : BIT_VECTOR := X"404ED56BC0CB88276A926C64DC5650001004745213082D740A0C165279B250D1";
constant m_0_3_A : BIT_VECTOR := X"000000000000000000000000000000000000000000000000001ECBA2601009C8";
constant m_0_3_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_4
constant m_0_4_0 : BIT_VECTOR := X"8D8143C6C04000A0820A0828A0504144014105140008A1012010014007FFFA51";
constant m_0_4_1 : BIT_VECTOR := X"089CC440890652131088080000A18E340A1E340071A050F1A0038C8143C64203";
constant m_0_4_2 : BIT_VECTOR := X"210856B5846DD32DBB0F09260000000061409240C04A0A0482024CA1210C2812";
constant m_0_4_3 : BIT_VECTOR := X"A1E0141822811E00490A0C40E84AD421E00490A0C40E8D2846B58C6B58D63085";
constant m_0_4_4 : BIT_VECTOR := X"0018D00031A03C018D00020D1AB0D86C3C23A1E00491A0C40E84780124283103";
constant m_0_4_5 : BIT_VECTOR := X"021000A250DD003C241E003A0031A000634000C680018D00031A000634000C68";
constant m_0_4_6 : BIT_VECTOR := X"424037045001284802020003A20C22000410171C08903890207160C70010A001";
constant m_0_4_7 : BIT_VECTOR := X"A4A000348902D6B58C6B5A521084294A524201A880028A006A28114202108A05";
constant m_0_4_8 : BIT_VECTOR := X"80FFC301FF8403401880180806100C000000D00014030800C00014000028000A";
constant m_0_4_9 : BIT_VECTOR := X"811304000D204281826002900081A12023A91685A01230169060804C010068E9";
constant m_0_4_A : BIT_VECTOR := X"000000000000000000000000000000000000000000000000000142588EA42216";
constant m_0_4_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_5
constant m_0_5_0 : BIT_VECTOR := X"8E912BC748A8209410894102944A08105128205140A894150924A32A27FFF815";
constant m_0_5_1 : BIT_VECTOR := X"020A111220A1080848A720F82095A634895E348531E44AF1E5698D912BC6CA69";
constant m_0_5_2 : BIT_VECTOR := X"631AD6B18C2128806000A8A91FFFD495532A8A10282A995440414295148A6551";
constant m_0_5_3 : BIT_VECTOR := X"50151B84664B015124992D049429309015124992D0494522C6B18D635AC6B5AC";
constant m_0_5_4 : BIT_VECTOR := X"80B8D10171A20C058D1040830628040202A25015124992D0494C05449264B412";
constant m_0_5_5 : BIT_VECTOR := X"42A10A892A128002A22501250171A202E34405C6880B8D10171A202E34405C68";
constant m_0_5_6 : BIT_VECTOR := X"2A081142CA8125010240E4A3082508C95452964552251A040A354A9701242894";
constant m_0_5_7 : BIT_VECTOR := X"806A2810AA42D2B4AD2308C230AD2B48421040AA2BCA59502965534A2B5298D1";
constant m_0_5_8 : BIT_VECTOR := X"BFFFC101FF9081040A141921024205048120440810832120D40830A290620419";
constant m_0_5_9 : BIT_VECTOR := X"1FE3FFFC7FFC47F1FFFF1FFE07E1FBFFFFFE0FFFC07D7E0FFFC180FE03873EBD";
constant m_0_5_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000001FC7F1FFFFC7F";
constant m_0_5_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_6
constant m_0_6_0 : BIT_VECTOR := X"8CDA49C6680AAD2590D2590A0692C8501A4B21504A81250400168A4827FFF859";
constant m_0_6_1 : BIT_VECTOR := X"0A02DDDA80A14B4B6A340082AD24AE36D24E368171F69271F54B8DDA49C6E84B";
constant m_0_6_2 : BIT_VECTOR := X"210AC6B58D764AB6ADA68081400004051A480A502220D2405311021010834901";
constant m_0_6_3 : BIT_VECTOR := X"94D0248526494D012499244526A55054D012499244524C084294A4214A521084";
constant m_0_6_4 : BIT_VECTOR := X"AA98DD5531BA95558DD552A54A0A45229A0494D012499244524D340492649114";
constant m_0_6_5 : BIT_VECTOR := X"40B982000864A49A028955495531BAAA637554C6EAA98DD5531BAAA637554C6E";
constant m_0_6_6 : BIT_VECTOR := X"486015509201494C025300232029A8004052965D52A52AA54A54081701B40C05";
constant m_0_6_7 : BIT_VECTOR := X"A6E02014AA50C6318C631AD6B58C6B5A535300A2A40012402849010022400816";
constant m_0_6_8 : BIT_VECTOR := X"3F00027E000401400880190806100D540500D02034012900402014028028100B";
constant m_0_6_9 : BIT_VECTOR := X"EF13F7E27DE27B89FBF89EF103F1FDFD37FF14DFB83E3F14DBE0F07F00004041";
constant m_0_6_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000001E2789FFDE27E";
constant m_0_6_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_7
constant m_0_7_0 : BIT_VECTOR := X"0081210040000890000900008048000401200000000090000000012000000001";
constant m_0_7_1 : BIT_VECTOR := X"000000000020414002000000089080040908042000204840200001812100C040";
constant m_0_7_2 : BIT_VECTOR := X"29484294A421201224A000204000100001200004000009000100000000002400";
constant m_0_7_3 : BIT_VECTOR := X"440112012601401000180440900014040100018040090D2A521084214A5294A5";
constant m_0_7_4 : BIT_VECTOR := X"202010404020850001041021428201008002440100018040090D004000601102";
constant m_0_7_5 : BIT_VECTOR := X"402902000212248000A440244040208080410100820201040402080804101008";
constant m_0_7_6 : BIT_VECTOR := X"20221110482124444201000B0000020000008604000008000010000701240800";
constant m_0_7_7 : BIT_VECTOR := X"A222021088125294A52948421084294A52111080040209042824010000000801";
constant m_0_7_8 : BIT_VECTOR := X"0000000000002341188108084210850025084122142109084122142084209108";
constant m_0_7_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_0
constant m_1_0_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_1
constant m_1_1_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_2
constant m_1_2_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_3
constant m_1_3_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_4
constant m_1_4_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_5
constant m_1_5_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_6
constant m_1_6_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_7
constant m_1_7_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";


end mem_content;

package body mem_content is

end mem_content;

